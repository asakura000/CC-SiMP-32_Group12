library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Common is
type processor_state is (S_INIT, S_IF, S_ID, S_EX, S_ME, S_WB, S_STOP); 
end Common;

package body Common is
 
end Common;
